--generate a possion-distributed random number, given a fixed lambda, when passed a uniformly distributed random number
